module tb;

endmodule; // tb
